`include "uvm_macros.svh"
`include "fifo_seq_item.sv"
`include "fifo_sequencer.sv"
`include "fifo_driver.sv"
`include "fifo_monitor.sv"
`include "fifo_agent.sv"
`include "fifo_scoreboard.sv"
`include "fifo_env.sv"
`include "fifo_base_sequence.sv"
`include "fifo_wr_sequence.sv"
`include "fifo_rd_sequence.sv"
`include "fifo_virtual_sequence.sv"
`include "fifo_base_test.sv"

package uvm_pkg;
  `include "uvm_pkg.svh"
endpackage